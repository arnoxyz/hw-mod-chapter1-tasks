library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity va_tb is
end entity;

architecture tb of va_tb is
begin
	--TODO: simulate vector adder
end architecture;
